module util

pub enum InputType {
	one_byte
	upper_u32
	upper_u64
	fraction
}
